module registro7 (iCLK, iRST_n, iENABLE, iSR, oPR, oSR);

	
	
	input iCLK, iRST_n, iENABLE, iSR;
	output reg [6:0] oPR;
	output oSR;
	
	always @ (posedge iCLK)
	
		begin
		
			if ( !iRST_n )
				begin
					oPR <= 0;							
				end
				
			else if ( iENABLE )
				begin
				
				
				
				
				end

			
			
			
		end
		
		
		
		
		
	
endmodule